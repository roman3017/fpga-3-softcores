/**
 * PLL configuration
 *
 * This Verilog module was generated automatically
 * using the icepll tool from the IceStorm project.
 * Use at your own risk.
 *
 * Given input frequency:        16.000 MHz
 * Requested output frequency:   42.000 MHz
 * Achieved output frequency:    42.000 MHz
 * out = ref * (DIVF + 1) / (2^DIVQ * (DIVR + 1))
 */

module ice_pll(
	input  clock_in,
	output clock_out,
	output locked
	);
`ifdef VERILATOR
assign clock_out = clock_in;
assign locked = 1'b1;
`else
SB_PLL40_CORE #(
		.FEEDBACK_PATH("SIMPLE"),
		.DIVR(4'b0000),		// DIVR =  0
		.DIVF(7'b101001),	// DIVF = 41
		.DIVQ(3'b100),		// DIVQ =  4
		.FILTER_RANGE(3'b001)	// FILTER_RANGE = 1
	) uut (
		.LOCK(locked),
		.RESETB(1'b1),
		.BYPASS(1'b0),
		.REFERENCECLK(clock_in),
		.PLLOUTCORE(clock_out)
		);
`endif
endmodule
